`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WVexAbNfD2ZsHkzzLLyMQZ6sMdA7JlAREWHyWmVUz6CFE4l+LzYQ6cToibtYQviY55dzeuvdHfmL
KDN7AJbD0w==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hnm8I1JRf67HZXF6FnJ/Cz4Fd9M1ehdX/DYLY8iC7j/bo9ylt1gdMWcbUcZiJ1De/go1CWd3w50U
fILJg0b8y/OjlL2iZbZVpLmIKwabWnzCOxTYCT7MRlQSScPJB5/Tqw1B2cKr68N+3RBc+hcxnU06
y1mbpmfL8LMtCwbQ5yA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f5TMU60DWU10v0OgxkC5bMqbLiuHP693vCWc7u7BXLcGmTUac0y/eMjHmNKM7GHjiFAYJiQnH8cB
W8k3H2Em0tQIOvYG+AauQQYxuy65ATH+VojFmw263AeadCOLijRTBtUknKqTyhqDORB/r4FvSwoh
faFqjbH/YHjNWa5dFexR//cDPrwQLUz5M8bWC2P4dLtosKwm4m8jGMZhfSS4WbQmXYISLbDZyPiq
y7o6KGbKmsqFzH67wyGhi3WbyaNMoJj+nVxyE4kDkGbJQVeELVIbj87/NPAFBpRwl6hlCOMrxaOz
TgH+Xu8Ft3i0hpKaPBpH5CGQ19hV0iJqrw7/Ow==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nwMpr1l4kKYa4PvrzMFQmnCIq9bOxwQlwrR1FnL4djwOnQxkK34OBX94Cq4CLIeIj1temHQ9rCTP
A3Di3wYCwhXTv3e3vEIYZS9SaPJnqsNmiLwmI9wqmXYdNM4xLA8UkM1AuPtPnf7IQpNor8v0t6c2
KhX3ZmtgPjAs69QB+KKVKbEOFZQ0Eo1J5pmjgKE9Wnu+RmgqgXNjDm9bqWeWBrJv3N71h19w2Su2
jG9eyMla9G8A6euM/dgeUD3QL4yCp5N7EY2n2z2FLJixRkrWV1LbS5kEH9jYjYVRF8zOMiVYNB8A
WikTIPaCwgiOwz5LrbgIgIWN72bE87LVrDj0cw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hj2NW6TzR3U6K13eowk6uRNnhfqMl2ClxqVmRoT59jmHME/KBizw7bRN+12db9vSDXcSCWPd2EXX
/rREpHORNh1eaJq46uU741+1ocgTt5xUreUjlppbtotGkRbmIOQ5sVvIZOhMQ/Z2ptGvAbxpZN4u
x+xrE5nnZj7/wqVPacM=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EXivfZIeZiK8X54eiLF/3M+S6Ps32iVEzFg2tGacWWuKBlWMhCgJutfLfZyjc9MnKjZidYa2Wi/Y
Bs0I3749s7dWdsslMx1Te+unGGe9mv2x6YvziIWON0/aNpP1o9XSRfW+Y7Wwm3K1QlFjswCpG7Sp
j1V8mDBGRf9KBJnTl3XBW42u8t8M60feqdsvJOX9xg295jSDUcd0kKSI4DVilOt1QKQSyTg9/7H6
PMBaPjPBTCWgkhXQlpPOosNDUDlmngWsZCOzvJ1mhfpdzSKszOVo8HqKYIRfzEa6PHzWwaHNJDHu
xECN7edzJtOJvvI11COLVdW5vmqy+mnLOtVuYA==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0UV3590fVcNIj9Su2uqMZ2sIHuEJpzucizkIJhzhY6ND0QDINgwc8A7XqRB+VVux+r/5ULMeOfke
dKw61dXzNPV3gyXdjBDqVDCK2jGvTVfyIIJno+1iWp8Bug4oWDEo+l0JJHdf+zzinPyB5fo0E67j
kPksFmA4nUh1RQBnNlgcvubBnWodLre5eSrvrPV06YZdOcZkNBesS8Pa8bjZqVcGSmoyvH0ia+kw
IJXKNN+T+5/UDzqVGoxTWu17huhRULRp8kqPPpmySPSzlhZTriVM+m2jfB3r7XptYNxmg8xM/ide
oHw/TLK1QEMexK9Lab8L6G+Gm08ixIz7IlC2YA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ieJJDUV9Y7y3szK6slyjnSJN5u9os7ryDdcWFwhmwPC9BFkjpIIIyxu9r7UTsw/pvOZh6bmeMiG2
W9809PpCtIovdu51b7rIsqsdbLh1za5z35aoeLHQ0VwT32aUM1Bxi5vuCDlSvIp6w1BAvtYYz6Ud
y88H4Rm2ly+Y6nQC1fbkI0mPo3Bp/pYjN2psvSELt10Pct3jCig09G/QpG09lP1Y57ESwzPTUH40
Z6vNivjW1Z+v7Os/U7NND0ZF+CZ6YFTdF8RiR3AWDc8Yo/88ZPjqQFADl+DS4wAWiYUwg4NhwRn1
/TkH7M59lKrRMs9wA/yl3ypR4I7dpdkUkWvZYQ==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l8PFcigsF210iXrFNZcc4DWio761YK7z4UCKqqd0CywHcwH0Frw7UgkCPg66symTJSlpO0qBNCJ5
/sbympyxpV+BwuY1x2aPLoOGduIvWJbE21kqRxtW4YyCLHWyh30c9myo6WJrypc6t3E9kPqSi998
9XAuKEV/VIKnYSUenMU+0IgAMy132UDFmxRkLrswTdPA0zy9Yxix0Tc3WXlcMqKuHZtjqwpXtDNA
3ZSXAaw7UERyMMPzDzQB3ILLivZJbdnqkYqRMeKi+zX4ltbkSufP7lOHa01ZwYMP2Mr0MJcDnY9A
msFjttobp5kjHO3SysGhXQ2mlvTLZ5CoxpRLeQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 28192)
`protect data_block
uAulWWE46CYoexUZMCTpEPl58Z3OeBNJLX0M25BizZr7wwR7ltVXNISo7dQRds3oZhbMi8WDrxgw
ptjO4+LSw9z0LpFH8sXv9sXoQ6kkbiOnXmmJZUaq2AQXMKDNZQ/DYDoVjaUSGHikRUMKKY6fLOv5
WSKk5dwe76gI9GdJ1iGHiRzYkZibPfEhHbbSqkG1UvIZ/Oku61O1DZ+F0MtGNct6fAj8LWJkGCPr
m4lYpw6DVxWGTyYGfnXVau9M7FO44wungC0u3DdwtklJiGaSW6chpsyw3ORa+JXtlQTAX+gIMUrI
K4Pu1xkxBXVIzXAHF5KoSTNBfrctNC6Q2VRM7RVu44e4BvDVhgW7/EVSxFxdZfCp8tM+PwHrokHy
A4oDEah4TKTsvJUiC4pEgxjbBQsLzQ5Ve1kIi+kis8xvoTQKqxGlxm2B38CK7izxFnWhR2acOiNK
i2cyV/82XbpX8xNPOtYuwZUxy58XIjXuG53hUePDa4BCZTCxgG+wC+uY+M/bkSS2ka7uNuYJZnxP
bPXTwxWF9x2t0H9hdhEBAhw3SfWouk8Bl1QE0oZBn2EhQZhb/4xQVE+1/jGZAdCxcW0kEPjjvUJG
K8VkEuKsKBiyBlwHVG70l6d5lcG0OxKDBH0sLmk5N4fAlqaa2XGZPHH1DEKPb6Pc6hMyFt0MpuC5
DLsA5DHjwtBP3i8Ygtl+b7ipVl4+KvPc2rgH0yB4LM3EpuzloQQvJC56AMVuytFB+ygWiJmDzmAG
n3KjPZCa8nAvZoUVPnweYYQPfcVc6tT42B+JWLRVtvWnRJ0SNZex4PYTfMhNQrO6p9oIyXznWIDZ
BAlMNNQem4g27k1g0lG4UOLvMKIE4TMTJ++RqLmxdPnfxbEsTNcGBjSuU5CUaiJjqAPDbKRPCT+k
tT3XT6cMnIn2Wbw8S6YMR63eI+LznlAjTEisMuBFUeqy5EK3BinAKELpdtY+6yt6YF19WfLJmjKP
bxVBZujTI7bWs4T+6+CB0fxsQcX9kOXKuBENseuXNpsSskKKJEGs0gifAsZDLEqo4VqtJvphXNgt
X7qpuLPo/FNSbw7kRxCZliTj6CUp9ICa5cB5XRMxdds/EQ0hMLYQCGem507sSYlxE3xHjIEe5V+C
hRRl7dH5Lo4BJHGszJpa++RKpHgTAIShygvaquecaQ1X+n7WevkukJVxSbDdIHVpN8dP8ZrY97Ul
rYJfCR3Qt3S1teaMAfaphjK23defZb5TNIE+KVQMP7la/rYC+ZY3j2JPZGojgYQf9/kPoNjE9fzs
ioBR/o89jTk7/ksSF2RXnt4kE08Mcyc1ZTdD6MjVKMWCNhTKtG+Ms9hh45eGlsRF7YFPUWTF3Bzp
NZzogOp0RY8eAehFFKhvkCOVqyurOvzb2jsbhehU+a/ZiJsemnvYykFMW3BJtAqL7kxgvDg83h5q
YXEaYhKs9gdIK/YgLcuZvddf8KIGJrqFMBx8fu1a2i/AyY028U+79Fi4JJwuvil2m2RjakJWyuaw
npFuyiZ8hf59Osy6Txs899mYODiUindExlVOlNAPwBHraEb0KeWT0pCVVfhd+g/99EC6eYSnv8JY
OAVAJj4J2q5Pqbl5uM3DQE7OuMOmwfNbpcBRxxuk9nZDMJtPDUhNGaq+sUs6i8IrpCtc6taRrCUc
QDutz6629ESXyZ/fdOkiUKxebb8CEKpwnOIDdXy1ENaUJhAabOXQz9vfe4Conj5bFSs4IWd3aMy8
Mg1Z2kA4j2bgby53rb4lYTYSVZvLA4ojVWk6LDQFkJdq7KRQWsUPOmjNPx2SHaAnhiZOOfArlzL3
hNTbgPkylcLC8hGMj5N+TqR6cdhmkB4UmpZYMwRVN0DwVqJLQbzQzL2x5NfDrhjbGFako7eLS2F6
LqKtrJdPF1Rz3eBvYcGTOfr/KQxnWcuKFbPZpYExXMM4AzS460HvCt/3rLzDMSQWXAZb3fdNLNSL
jBqhBDAq35YMj3G15tabJUjKEcqqrDX8A2FMhqa0ilfOm+R5BcEUN6jvEKmNHlYUysRqBG/LgB4Z
0FMLibQn4br7G1kW753Vpd/BPVmGtCtt8t8XvLiZjaJu5hQU+NAF+tSgYB7OkfoNb54Axb77+2RU
AUAruCTBoDNfsrGFzXeSnAOLN+bJGdZ88xTxLhE+NOHpnewbgvda813O+2pmY88ECWBqcz0dphbz
uklC/mJZ9Pu4mhyNYnfqx75lefDlALhBMWlWaWz2YMzENlyqc9Br98HltuEzgVY/1Gzq+1pqSs6C
vzKVHAwnAzsqYGG7Ed3+HJ8sOYvFHUj+5ay12YlHGGwO6zO3/r4c3vzAWVg3v4ips+pBCP+orZqs
QtNMQYkRAuPpUl6yA2ZvOgAtCXf9wqEb+sCPBSwe2Ix7AlmTvv9OKSyZGYfEssr8X1vfY/IwDuaY
QjbaKwM5F+pnklTvI/L4Tyj+aVVfNZAtIrcLZv3kb0yUb82Fa/nKvGSoPrB5oks2Hz78gL3nLuaT
UKqRlK59H+9JFAgLSP12qX70lQ69xD7QzHM1zS3GwQvgVpygPJNFt5ihBEhuPKr7/tSuQHkfmBoE
RL2/eY6mFMpw7kXmG8XjHp4rJlu3d8NvfEa4oDYJGj30LC7oEnHy3RYsoTj2gu2PKUOQmXTsoBDa
t8XXeYRIBrRuuIefw6Lbr1b8Cxk87P9ucXPjisNLCn6TNsLGhnDr3To+eGOcdqO2Jdhhnr4chu5O
E82WlCbhcP/GUSr1HlNpOYUQqhdOS+5YB0pP3358bXwjQQIuhEYN2UEwDGf2fyI41dupumgRpsMV
pLU2/AXtBOT1obFBDWtKQcEriMoW71KXG0P3228b1uPWxsYDtQvK55UYpRVP19r7g/GHcEz6tvhI
vAVEDpkMe+08ZHsDNC3KvvLwaI9L0y1XVeCIoXEyNKYXIW1OLIj+/hcs8gEXtBrNEG6uuzE5/yib
i1jdSc89twhkAulMbNKevweY/O6Z2i2oJsWORJI15QZQSvC7PiDkKxG5mLtMHocTgUZmJVw8MoDg
mNJGTna+q2nQQR5D9IWfGHJqxevDzo/2DmDlHsVND6awexqCkwhvse92wvrY+xDIs+NSZsylxW1T
WilWAYu/y8klq+A/vs415C4HAT81YdW6jY3M5w202fYovSypfP+nnjjbDih+tQwg2jhPlzHLFR8r
XjDV5wCKIeMqHdYeBxrbfvkroNeN19iYc8hNI38iJlsLx3Q932YziL4x27kplENxWd6Yn+lL90ec
1/wTsPjWMIv/+Y5kxwCk2H1ET1+yB7/Hd6cwhhvDqD7rLAYEORltkgaCweEi6HuUlVkrOeLQYpv2
ljjrpc0NQIX3SjVzQ+YBlflupjmM5TsENH/bGOEL5zdy+1fiiWClruRqqbF+/rBFsDfZ3bzH+yVf
Epj2dlOVO8TsXfKU3BMgPR97wNMbOTzsOdJGOXhEvdCAw2YZQXOhuIV3nguVKpDTBdtzdE/zMzF4
3D0eggwShifhB/Q46SgM93v4xyPk3nElp3aMcDy9IIOg7n5mRkYD7RPYcXJ5il63glLY2kWFLeYn
5etPYiKrX1seM254gM/5Dzz3lPyMvUz5U7/Wtq+m8KfKsHNzgntFvG+dwsrAI19twSTOAUkFj0yJ
ZpSfgQZkpkKBNaAIW4ecMtFnBAqeAXTSNmZ3W5Yj94I0yhQs91HuWn1EOgyCU511pBsukgN23Gcu
hIcQ+IJbd+AYpy+0LlWqmmtrtxJdVojWuFUL+3lV8GgozAGBXGOOyANpJSXpI94DN5Yv3tVhDynW
Ez6a6+qqq1mFYyQIo/VRSVpM+ns0na0tBDmPztzDnqH439k2tpgmFEYaEHpEp0p3fygvegaG0Hie
bnxT0uI6mH+2KOxnGqRAunE/eTeu4qr6VvM3yWbZX9H014+876bhMzHP4tkY/kgic+NA2vIVdnZu
AJFQ81zjDhchvdjxcXQMoPlr5T9kuuJ/RaYp/9Vbn5VZ6nuFCQ9SvDhPmCk/ryCHUzv8VxTKzj2S
UXqgUZzZT20BQ4uEAnpQgmlxihttxJvl8tcrjjPQTXIhBQsaiXaxd5M1l+eI+FhzoXD/+7F5SQI5
sYKFHI8yH/4zIfMayLUkpSmGnzx/wjCQgDWNpHVY+A1EnFr5RfT/fAkYeB8cwmsL+XvjV9BDNgwE
K9+vomlglkuVWYUzzpR5vmKez6E7dO2J8NH9dvy8OjlpWQf9AWYva2dbyH0Vw5Weo36pCQL9D/N7
QFjyiao4qwvlJUXC0HLRZ2miYqOYWzAuUk/15gI2J4w34lmbyUd6BY5IumGp3fpCTNUNR3qfuHCj
lU28pX+vwdYyOX6DMeN+Vsv48U2NTOnoIrhV+JKv+rJlhEisggYwNUTZaUNq3xYuK1jL+ubt/W1R
LAe5JkGjW0wvZqbEp7gEH9TVIHq3UFDI7JxRS9l3l69+Rne+8r8MDN0QE9ILh87lnY5RmJrRQf/1
vLryq3GhG+Lfzb0hULR5s5624lOGOWFNGupNTqas574IwYll5QnuKwO9geJIDUBzOg1TTgGwma1j
cZwowZN2Vl2vELRQkQgOgL97wu0oI+La437Il+0kwYhMcRmEly0wrZfcohYTx87XlciOAPlpj1zN
PtirDA4JrMdaIicqVNh9bUaFbCLuUgfwcc02yd5ugOzmTksJZIYtbKD8rBZSnzO61S23mbEmShvx
rlW9NxtngyoAPJ8OB1lLl3GvZonTKGGXJKGppqyXr79CLUmOFbR1z+Beza9oAkgeTfdgSTYTlP/W
wMlVaphs3FBuLKjMsLkmh17aXzzZllUC95UtN/GoZyAKNnQd4T08FfVzEIo4pGneTXU+1FAj/SPw
JS8mpZAMu03Kjg5jcg1w0iyy+2BUdPo6vsqcTsWt87ZCUonh94vqyfQpEPn0Snuq4t44epRWJ6a5
mxs41FCDhH9zGXUO+nM5s+rUh1DRSrasFFiU4ZSBQWbOx+kBLDqvrYm7itm7CqcaBAgDlLLeg8MP
rBGBYzuEPeKqwzcidULuihohY9ioxwAW2XuXcaHTSIkx3iqhOQ67PrIbbkw38JZOheOX4t6A3d+t
1ChhOqKxDRGKexIpOs3Dc80bFPIyq6fGVVIS5Q310uVTGKaXeV/qw/8+tYyu4EbDQMhSiSRL0CuQ
/mbzFU4gcG7tJBEC70bv9D8XT48A0Y76nXAJTZr8jXQnEbUNGs24uM3zAh/SPV+p+HrfaI7kqu9B
aSPJE+EfFfnGtI1WHZ8iw9xxV7g+PedYl+y8RuHZmJS/1vAu8+y6hVz7hzEKJ3yWfSIQp+4+5pv7
MriFqMfD25sw1EzAufat6lJUwHKY74c4plFYDRpaM117aBJw9arTjwhHmjDwQxzxOlQA2OJ6iEvp
VXJv6LElFK+vbWm1nBnBQvXqA+/1vMdHFa5jD+tRqCrngGukGcND/ZnVqyuQGU158L7DtcbbE5wG
gNUYKX5uYMpLdcqD3zsWa81IBRrlUcs6a74n0uDGwagdnq3HAJLvpHx3goPIfLiMW94raNzSMunQ
3kvN4hqXQpJFAOKg3nDyLK7CY/Z6XgBurDCW/9EmzAE73MK7dYACHzIJCWy7al9bT5e1DlfUb+cR
4bEKrR2KI4EySxR+3sv4gYF8MDNMgHvlbCbDOrwe03XqRxbc1RWk2/j5R/jEcu1nvPCkx0rmDHZ5
rOOtp/VEiFhuYFVuRRPhO0Wgq4CJjB8EwwvHY1eiLyKxP+j3+LqNXcpuzazSYKWd5vhqrSFLQuik
Q5NJeja7ExdutCd/+5XoXNw3PelGc9ZAXmkk0YLb/jz80RybSiegnA39/HG9TKS2qk86ziV4H0Yj
KoyDRKVC0SUaGoqVgMy8tNwVVeyh+Wlk34WHjvri7RwxkHuLrP0JZ5cxFjPaZxCumxIscdlPCt29
pv6P+XbnVkVXkR+XBIBwFEpsP01mlq5F1arP3fGYT23kI3WZFy+K7JGABadpvwf1IwDTh9BM0rqu
ICqHDoplRjS9fA9P3r6vNjReEnzSfcurH6HG6UIhsjcUJgskE2RwV50SirQp9KImjybp8yX/DkUi
zYitNYQvjnL8kjhswUE/2IzwLG/812/Wo3CfyFS16671l+Pwbtwnci7+Q3cvOMHv5kF4RIoZ/XS5
FQOJe+z0JtPd90ZwKvQU7a7g/Fo5YC/WUFL1G103BwKYOBdUEdO/oIqYDpodFk2xX1qgk56TiwPR
6T2GVDxIdLJ/9kII9XbznrPVTanzAwVFZoLrx1v46R2dyJSrmOjQ7Vb9IPyyeDukgXAXDJfmHAz2
GcytEHiBf3tx6DYTpTBMHCJWKKuRDdcRZUCCOZjh0Eyb5jViaFHCAKr/+PUUpWFNyjntzB7GS9A+
HW5RBbFNSANReyVeEJukfXHRG1t1Q+s7AAzfqkx0JPCMHUgtiw4TpMiSn1rXRTX085RN0gvvYPsu
LkQ1ILJJVdg9dmTGSxghGYxSmlh30iHNbYwrG1IFYDFa/DfBUAFNWueQU4+i2z2o5adgiM4JJ9of
1V+HVUA8ADCct3mb5enptJqG/Sva5YpPzS+QNKA6zAXllvw8RUuBacqKkgcMaQwzev51cd9lNka4
AxcpQ54AYnEsIvE5GEHTzG/9G8TlZcKXjEm/4kbZ2udjfJ/0xVchPNjaOtg5N1Zs/aUN/5U6dpJB
G+ZJjgmZCJT33DLMZNI5ImpvNinW/vDyrkiG/1WZefLYpzJeXxN/wtHA6yrqelowHpy4c8iQ5ye6
QjxMwbY/pkMToaIBIW2ha0PWd4FEczXam7VGsZTubVGxN3RDK00D+f66YhMD3FfmA+TPdDbvI2Rs
Aa513pvoOa3Mp/O6Lf2OacKIYoVs9kQSB6PTf2kXVwoLCnHdY58Te4MRfwD1jUyH07pCWooH48XH
aOm9ByL2exgX73axf7v89t5CQY8/juCu7enFaNlf6bNC2I4grhb99/qyJ5ybhCOrtBZsAM0cNjqS
H+z3Np8L89GPs62gLMJXj8kXUqupYtsom30sou+WLmnc5b1+5v/i6RWDU6++sWarPljWn0UYvtil
qB77EkIoByS6sEReREW7PKSTWiuKMcO7CMRDqKY/4ugLj+KaAXtte8Q+G4rSBivAG7UX13M7AlQ5
MylmUp8A8TiWLVbr0x8p0lZ4qaEIkGx+gKCSo8A9ej6DPrHiLfhBdjWJKsu9BCaXy7KeWu6rpnyb
Yyl+avZ0ZngfSLQkQ5B26lga7z/TBC76k460xWeoxPRrLWXBBxRlHNgmZqYBxNnTwXzkjvRvMcvk
Bi413zNuTGg3M+0eyGv1K2fhgKu7TA2SljLE2Mq/levflKrazvQnxMKR0qYoPX6PShu6P7H+K5Cv
MFjimjGsG9MDe5oTvsvzNPDBSGgqPlO6csB9TCuqr4fwduTipVKXifyoreDAANuAQGQW5qPMVPnW
y9/VUi8w2S8y7aa7sNf1eqm2BsCLShQMPAjqwv3vOZd/hHaz80eIE7GsNb7mjUe29ASeduoYKPuy
Woe3Bkq5/j+a3yrynRaLqvk9DviA1o3PYYRiT4T0RXLW0glI3RUEZ4zob1o0FmZbBmDtmzQ0hXLM
J5RiW8pftD8X99+I7GXlbv/MWs0/tZIS/0/rZ36I+RyMRVI8aYRFkCPD6iseEcu1aH3STOaYyCpo
6xHdPzlegxYRtgBiJsGo7q0zK7YzEcPrc2XiEdBowlk38m74yAzcTtkwVRIffWYppT0YVjuDiy6E
dYRCGaKdXZj79tVgGgBgwKcNTQ/wTBnAak8o34/zeGow0+Bw/cG6OOS/5NK4njnLO8Ajly61IoBD
Hj6dy3jFXgA1ZsBVZbAgOlzY7QaoEdVSz4UXV/zwKYQzYtzLc5+QBbecau3FLILZZkKFdndTBJo3
OO+UxtsdHDOg1hA9PMqlrNitmDDIjZ4nVyVVbje+xBLStqd69rMPaSr04UV+PS/rV1sx56bFFvoy
fbZGjbF56KkByDyg1UdcZfhGV7xLXCagdts/YVIptb19Uw/xHPp/oMbAgFOhrojR5xWr5bqObv+t
s/PrkwQ+d58T8cF70L0xoVqwKKzJtLckbWhyjbYZF2RuOd31EpvQ8FgCRYlEvcbx0xhgkCgmKm3G
bEFe+/A34QCNta4BMQbhRCiuSFtEoEbqOsXeufuxjBi38Zimlchcti/0Y0w6g/bI2L9IeGeSwG5T
k+7J8SiV9QMRL2TLntxV+p7w5jQH7N7fbdpq6iX8QkrudSz3yxNxqUAdmyRMi0yQoh0p2i+l33RP
otV/chFjKwCBSRwXlkDO7L0bI9EkfMhDzHBxghZiHcQc7voxS4W25h+VsdZjFmI/sX/dTubnki1M
U3ZVSHL1bULJ8I9tuLqlPuHCUN5it3m/0ZYZ4lfQdyVSw2Ah8OH6/4YNIozbbmxGVQBO3EL4AFxD
ikqowwYgHwkHBBcbB9WG++KCL8kNjaYLPAFfJ6tIiRi5xpMGYmnfLpuaQ8Vjzv6HBtGDu1lm8Ais
oKUanmG0oG8JMaNyjsFgDYQfjOC5VFhOcCnOflGpiuSsGu0bX6bM2MyKwjgMAQi8gpY0qeu2DF1a
qJrygwhT0J8aaf2FoY4IbCzhA9xMVFeoc2Bq1MX3ZoFJaynfXEw3IzB6oC95y5TAN9dKDY4DWZU2
0CpWcqLgJQwTZyLd+iAqkZOeeSv9CRS3ZXW64ufvBaTUtvqEcj3j88U12vgX/LWowRA0ND3h1j60
m6SbOwLxmv6kiFdZttdiNYZ05NNeswILr75jE6Yi3GsKZGGIG7duR8xrwMMkfHMZ09ODcC6l76F5
dnUC3m8vsmGZ2K/5ViPatDp/xdF0yZcellSprWDF/F59v+ighCtmN8vbe44Q7CgApzvbphj1dc7J
guM9i5DoNjoezmexhutEAknmgYyW3+wFqdZCFPVCZDBTbbQrd3wafvqxF2OcvWNmKm3trhjmlIKL
ylREsjpL+LiOSMe0gHULffJhxEgPEuWPF9LQyItj3VdjZ3irE3amwCatKWB2Q/fzLtJ+W7ynmGxV
l7I8Jgbfq5mGcyytYegCaCB6iwVlLoXLdmwCEDkUfhDfQVmG1+ZrcW3OlFtNT8BniDeHpAzkS/Cw
SMRmSWRinX9zX4pW0NzRWVzJAAHsUYyvBrsH3ANLdI1VcSdcqaYW+ifcp+ujOfKpgLbBdbGTfd3U
S8K7A4IpX5qbzl6ndcQu0u7VKOzSRpFL5pFZSfochCnktKxfodAbxUDLND/hQqfz9Ybc4nA/ghjg
ZBtvcxIbjrftiCQK98jX33FqcyoSAd/nWrdiRvmYUPHufQ3vKiXLcUU5VP+aZbetaW6YXuSF6RB1
2WNE+mp8mjz8l2cyY2mhVlrjft0/d6mNW+UgoqRFTBjbhcD8tBFqOnggX4rWvN01lccFwXBuXtr/
p1dLlQaKWPOrEHM0nKCyjl7wLAreSoJlLapmB6dCX91tGoRZt5Z6KMBolyA3AiaW3/ePQKgfczs/
WgezZTirrVit5bZ8iwY16PAG/6KQHmv/kbXbkggzzicXjgky2ZXTi5g9RgNY1XzI2B998uOdlq+u
4hpB1HEh+no64lnk6RZbsz2sgXCCov0ny1khS7vPgSn5jpaWkPIwYImgVDlwuBO8GBbDd8+hPs9j
CJ1Jf5kaoffhNgUqyuRCdOTk4bbGGOD4QEia6REKm0mHXktWt0eigdeJ8GZWJe3dCpL93ebyfI+F
F1+xrLQUD16Arv5s9pZwle1fduQjMuOzI4P3X3HlfzpM0ncnVEVA685LIgOnB3v9KMBZ/gObZhWc
RlY8DjiqidGO5+5VQuHafuXwy5EmDxqR1ZySG9RYoliEogYTetU2Nrcfc4deUWiOZ2917xi7opaD
UZS/JjHdUBAtguKxd3FFn+adLbi+3lJ9GrgQHgKp0TF1207UEDGcB1h5nMWfy3HLueN/Cit1+4MQ
ZhvidW+SOWk4FgSXcpk16kHAuZ6tjogRuMEuhpwVfZ6R+gyaEGCYRba5u+C18yNXZfLTEYo1x+Bq
GNxVnLPBbwXLot5MLqMm2oqYxSzgNBhMoX233Ose4X4O1w4cOpg3KPeLYy8LpW5sVf4Pgh1gdBQ1
ikUVkgSJb2P6Ty6CfNHF7RmZwfG6WHA+aDkEj6N66BenyvEK6U6yFdfESmlTZkhKq+Zcfrd2ms1D
bbbg1UMBW9NxUrs9y3g68koGdv/6yPFm/nusbjfSV6tzf2O+V01iT+WALrDQFDW9f/VwNyf1Qb6o
H989XJxqcyZyA7g18A61vVSv8BrAWDWymRvJtPa44mXRbZsNAJso61WxqtlRays9IuCcisVF3uMc
FwreyD+mgo1siI32F+1kvNFMBwuvVECV9TpcSegbhkwgWy9XXRzDLT6n8KyNZbBzDIFA/2ADkpH3
NzXEGzOJQBkx24Eihoi0r/ltNvHtODsY5b9BsgAw07ZrXUJTeYXamwrett2u/73yrC1XDenlSi02
c3YvmfqpLyzxPXZLoUv9nuz8YzAttvn0fJ9Bes3RgKDVO4iyFPksz6H8vjG0Kg2p3QcmWWhBTMJ0
Qncj1yxnGQu016VhakNyYNP5UraxGoh+JPyptgbrb8hgymXaX6vh5JLP8fNusCjV/MIQDy7jPZ9q
Wp+lqGu4PIXniAHuXI1+/ksIDKVHQnKgFTdWV4u4X6JBqavTo29OqTPRT/XSPqq7FtWnfP8GzUm/
b9Ps6Yk0Avbloq+XNNbPm6nxX+hhE5ExyMqtiSByWWNAF7qhknpv4nZlKTfyfdO5arNb3s20H1TC
XrWsXlnUw6cx3cT7T3F8mxacA3JkDcl+PI9XWQeHQXfVsxbKEdCjQmVoObo7FxUi2gTH19qbO37M
8Vzu7SHGpVOzTYtr3SACluXpHZ7tH7ZHDCSGcCi/an1vmaicsQmtryPuhNh6N4dD8gqfsXnI/7o3
j5shY/phDNbvBAsNoW+HDowgAJ+uFiBpIARq+Ae+L5waTESJ9PdJsg8+vfgcliTogcWANdxaklTU
MDFL23BWV0A8+JJkce+QeNwam61wbHndDsn0ksG5dsrt3WUukHXz+I5Lt0KwWaDlRCLt4KpP0L4x
azUp5Gjg6QyKhaJSsdH+bzKJ5YByxSKsimhplZuNCRpzLUr/utp73uNLztTMbpjDa5Vk9oWYbaWl
5VBoPla0VtouNiBg2qHecNejyrz5SW741Y4iXj2w8Y/tUz8mAmFjfqP5UVfywxdAjDzVAuaWmw25
4r22P1S+A5Pd1+TGnC2/EqtyJBqMajI4nZDqMAA+xygq40goAWIhgLQQEby3rjRfl8gJ+Dxd6OzL
kf1zckgt/KwRlfzF2rSyftWPzCpuae8d9Tga1J7eLuoNQUQO6MLTxNKc4pM3fwo7kVPRnAgXpnUG
eze4uEVSi/bI0yxqi70UqRCwTEgu+yxihGMo0LRmPRZLyNrPrMums6iYXBeO72IGx+Hatxerb/I2
g/hEIqAnKQRUcsflCPx6MfHX9Cp8I3dL7QaxJ2HmhPBtL0+1znKJl6CALTKQsqM9kRc/noF309Bq
LCSjoFwRvOn9c10Sumu4q+vC5OLmYfM/qkU6JYgwrHz11uDorRTXAq+zqlDhFKmrcerHKK7wip15
uYhv0oRxEiROTw/lqkIKT7j1tVUg5B4Na0sH9Bwua1yCs49DJzvhdd79pHS8VNq5YzJUN+uErgkZ
g+BOXmXruG5Rh2QJSjP+wTl+dNeiao0WHDPoyGP/PU1vFXVPeNPXM00786vrA7dRYHtB9qEbxYa4
bFAqvIrXRdWN1SqCUiBfz5l9qrNPRVvoUp4HiwXmbzK8p8RxgyDVqxE0w9FkwsQ1P65/qxOF6yL3
+AiDtDs3btM/XFkXVrZew13+jJLlRmefibUmHkVfZOljRu7ygbLpXAxwQ8L1gMn/h/7xveI7Npta
RMdO+/JXle3uU44xl20KZe2omJ8uL59l9bLNycvTcZhPVvHju7OK3itoXa9rJm9OT9998WnKyYrZ
j30i6QaQN93/UlqvUFPcAqgVEVwYSLNuWgIDsbpVJs5UmkBantFd+++gzXqDH8FvCQB3nbs90Qge
I+OXeLv71L99cs+i5q6yNLh5HZNUgx3Gx80zoD1kZYLlaIaUsTMH34cTKWKDoIN9dTgjiYxV5FII
fZYMZBTLHee5wY7pKcjOXxQ6bleWlD1a8FPWFW9a9pRX8D6pbB4IDBFFVetPgrCKw4kCrGgqzXs8
btuvXLUZdltdotbqa027EpACCiHnwA9i5fnw3k3rIaIl+BOnnWB2PdLDYaliq+jyxhG675y5skOV
xouEy5TnKMAIqluOtZKHyKa7fbtw8T/6Ojm6ZjZ2zGU9FLayU1GHDwAjUYInueWn/KmfHjSvJXXI
2kfzILbwsw4QhQz2VMXyJJMDVi3MLR+nnq28Vk4yPWs8nhRpBySxnBVEuuRWQN608tR5pIh4UXZM
9M+LA8PSQodYDXCRt9i6ybbwNF46B0WkoyxR7+eMa1OTWuTwNJRCTjc+KlclBNS9h5f6/n9jqGPs
1olh/aujMneqnUZY0bEfF9aRTyNGNQakeq49hQ+sdxzPsdRQSkD9nVvZpO48r/k/uFV1DreC1azP
jFdKI2K2hP2FwKKPl+5B2JFPtXMY6/pFL8acsDrj5mJ0Vw+K8ReBWi1ITdqub3V7iAMVQEv1pT4R
Ve2Nzoed2h0IOs6h4Gu7ptUR57WUfbuqEMySTfeL3FZrcYaCvd034B8x7ZE6B4b5JmJ9tq5zz0HU
HHBR8JqJ8WWSHL9aWUNmUpkCmmYfGtmgYBHXIrsWc0mHa12TsmnxQaZauOHnvxPtkxr7gwjYAPr1
Pae10NIcPuSYqoXeSt59ywC0R8Qi6JYMPH2fZNxSXaWmS9tpfMTmqTLUx/hHPlA/18P58tm0MiA7
gc36jERLxKwiXa2ZWUKZp7r+vcLHTHxpXpEOQbGH/u4H/QW/14DwfV1gHZttCQqNkTT8ZrQW0UNm
jfKdKnJ3UnFUIzrNWxcZhL5R7f0s1TMDxDC8ZfNE2Y8vNEfgJdZXwNMW56mMmcXtCBktNldGzhga
kTqixppZCaa23MY4LeCY8v0G7D682yHretqbXlJdxKPJZk3tSod/aV/4tjIwCTS7d3hlsnbl6QgH
ZhA7/uWPRt28t/5mzxa6yTxLG2I3ZedxwPpTYsmLJeqMh8SB379/Wa8Ixbd10mvfGHTvmXuPK8Ym
SMYJFEgn8+SQo8orJUfqHAS3i7f1ISe7A6s9TIJby5exLVflS+mT5pLRdQDhFWG762wrncq2AXOV
6buT9ougR4SQP41YDiyg8QhV/1/S8qqIa549PLlCkNPZ3T4EIuHnhUJzu/J5IRPo23Gqm7FpnupQ
vVn2Q/5saTwtzVKm5OGemfXsotVAeh1Ut3QebS0qJMDOidM/poK/kfazJnmnVHUhKPQg3g7umeFT
gi257OVqdq6VjA8yk0ELr71xp44ty2pdgLRbYz+xGXRPuqTqhDLA5eew8GVd/watR9oMkw5uZQFo
MBIrQxEmYARmvIJ/tb0vQzN2j7lD1BATdqbQu7sjpI0eJfHVntVBKBJX+Cn7DNTfN5OhPQbQUXa8
mzgLMkpgEc349Kf83D0ct05yg2sy+5yTEvt8QtstZrWLdorhGGRL8PCijvdnp9lMEBJ1yeJaUE29
cDydPss3E5OG0y85HgqduRWDAtAD9zsBIXzgpjjibz7hW9aF2TyV3z1pR2j7X9a5/SdfemMCvl0M
lAMToHjSbUBHZCH0WjaOpVpPRxQogGjyG2pyJ+0rhZNJJUFVmmlxEWyB580sp7PxXbvDUcwzuwfD
1ufBy5+c7utnaToqDg4jhh14WcR4QGmiBNojFwG06R5LNLPrGjrpNvXSKdqUe6ox7Ax46m7q4w6D
XJ1BfjlViY1o6vhN9hoZP10D3zBRSPzt64kZ7IHHLm5jmeJRi6ho/YlOx6G976dP34tfhvk6zFjC
rl52dEQizwoTf1ztkQ8/mqdKza16R87icLoUIoQ/pYQKb0nhslHTQfc16r6HJqSYm5vc5UwqGfxF
2jg4l6vzUQ1wIsNVAtpeUyNnZCMHpn4QGQEG82y3Q0vlS+LtQEA/ZYveqbBnK9VwMmG+y90HP4Z1
kG1nQYKGy4jiTqieblJ5/KQF3OiuVU2KC4nXPFt2soaClvn3AZn6a2Ds82xjN+onVLLyODxkSkY5
ew7/i0CpVSyjzRsW2Etle+aVtxCXTl2Mstl0pgH2582SCfRqxJMN9YrHPo+3b+/gRqopm5ejrkFU
MhNQ+DYStUxJJQu+kbPQoyVTpJtWsoLO96qeHwkO7Xdl5Z6CG/tOLSy4xuTfZYcRbKhgtTBcWWNg
urRXWD11WmXwLnt6HD2NobgTEzs1JmwNTIkgcqds0yfd9VrziwFcXTdDC8fUhWUp7HFDm1qcrN6p
sZiI5+d0dBg3qEe9d1EnrfQ+hLt83funCTx55dQAFVAFwYRj8xhvCCFRHHfnto1Kmu89o2ez9TsU
o/acl5vWinpw0vAI1q/M23KQocwByaNa0BV9NA5+K3ky02Ziqq1EjOP0u3zWBQwz2NvpUIxKnBK9
1VQXnqrE9FKRbkckuGqkhS8tTOv9148X0A7A37hXuEhivu8BczY8S0i/xm6dh3jCTUF/3rMytBUL
fh0zhQCNupNI2y0VBEzzKC07GzUQuq1HxL7xeUpSYRt6SYNp+7PO7OaZcUD0KEQXK3/jTQ+r49c2
jmhA3k/Eigncr34LiCMCdbGNIzbFjvigpc2xL7fzl2fTb4eJJKiWhLpGNITmnnqRw9cMHYmYZKZM
H4o6uCldop1BH2lFLchQ6XsYFL2m5HamNg8loIEUHjMvoXcn0hPqocUA9DJsexRSPHwuEv0jYCvu
IgnED7kD0mQBkhOSryMgM8xtwHQhPBRd56oqTSpOHMbnUDQ5PKMLcAW9uB/jClcKiDBAgTLz0oc0
3alQ5DEhhZoDGoR2IVIeVENdtA2lGYXfzKCB6XwoEsLtvKpbt9gPs+1VtNYtOC0gyO4tLsJ8PHPJ
bek92dnqlcpZHhvv7oUosteRkVgYcxle4qUL/Q1I2zQeCW+gi6QLEyclAYfltmufdrgxvjAsHdOX
1a+zy4shOGsc+2CFQhZPxGU4FR6eaTHyt/g2/TaUKDtX2S1LBhlMSsT/eQJaq9yRqzmMIRJJrJM6
jDkefmfmD1UovaEQjuPzS1XKnwqJ0AdMc9VK1a26HpSQdINiIac4D/w1QxgBqJrJihStasBlwKWF
fvIZ1N1Z4eW0IPnLUXXtGIHD0qF5R4CPXPpy/QIlE92KXKD4VNgBrxThbVq6iA6mK6Tjjh21f6or
MaoLeUqyqpklHDo9xKlbn43lARz4DyojncKx8NabtywRO7EB1Nq4MXQ+7ifsLWMU6vphvrqLKd/r
jeRRBasTwkt6qN7+CPett8Q0Wqd4WDhjNAraAZnDDumuMU8IJ5dgCZl58zAZcmte2HDB6YfdWeBY
zHvfoltekZqm8TuGnQw74AA1Une9V4XQOeNiVG4qCVLLMktA4m3nexj9T5A7PKwreymDzK/54umv
/5WibLFWNPQMjNr74FbKU3cuLKZIp2L5+dsRmm7Y7Bb9D1WINgFnk9yyKdMklt8DrOuTX2XUvAuN
1AKx6Sy5a9inBdLq+/gjJoHDPtbCwkmsUW/4p4A9oWRRQqXVjheIclz+7z2h4tSIySKRzzb1h+E8
a33Ivsc2p5qMl2dsca0SSNsL/GWJruAxTTiVH/4fzOCIwQMzu4MKidsxvG6FX8waU5VE77s5Y9JG
apxeH9UBIjAMbunLEv6/hkESwc4E8+ykuMdrYMq21sjMAiXq8r1+bbD3JR4JupVZhtXXnJXpGhh9
cAHp5u7O2Qxn6JAmbFR7ba0/l6Xm4MudiZwnLL6tL1sj2lI9//CUdbV6Ad9ELyxWnXN+F+7QPlf7
B4ni3wC54yC7ojmzYnZ4J7XhUKOcOiY+oZUEqiqeKO87ATf5mM8x79g4Fm4HqjRfoKkYmWVdPdtv
jVdevpnsPGt80ArTLwFNAv8HEUYOicw2IvOQ0OlGfnmsw4OA0+Q775slQ3Ll9feyG7GwxQu3XgSG
bIcwIeB5mVCeafzXFxjiY8sc+2xb68xjwMFIkAWMte04LugvVzB5LVR7qeDfFe2F5r20omi20hff
p9RkIwbO3WCvpp6Gkuo1XmeD5UZgc1syCDdzDBaw6p7G9PIz49keEZwwf9mWyickRNundqktJt/T
b6i1wx0yjGafEKutEkVf3Vs5Joz4qPp7Cp8yc2l0gf6fXqaA0beBGkO1rLdLD6z09apZF0EuY4ye
lN8YzsJGEeCsGWWvKAjNdkqVLBaZC/5KuqT/QhwQMXc2FiTe32nAesBmp6W+W6suKsCPfDsDI9Tj
YFCzXy2UvUq1JhXY54Yk6cwHRfnotPczVKL347FSP7defhjy0MGbu5XVeLnDRIYy2/RJMnrBBc6O
y4DfJW9LS36Fl9DPQ9M4vfIo77BIBQROUJiPB8De1BrU96a+HaDaJAGEw2nAaCx3vn5AEhxU8sAk
iEbstNJaQuS0xgHz7U7QkfCGqqoPdFlUvbwjm+xycW3LdQhCTjGVBABB1D6tFqG7vMF9GMFrw7Zk
BQSARbVPp1Esvd1CPKwo/jzGXDsw1q17Z3NCHsPrRZMRcpnJ8ZiLA4elFJR/eNZZR3ZSzix4Opbx
bXf3k5CUYCIMxJ8Rv+mw6REyIwGQG5jBvJMLWjVrJeSHkPL8SjkeSQSa+gonjND+kxRXtoZNlP7p
o0DLBUAhYHR54x4UZZLOBxXdtv2WoZ+UXvO54w3MofJ+x2H91ju++YaPOGJI7uPXkkysv71u7Uex
XIdQm/YBzHFfystVJGW02rF0hu9dWQ4gjccSacqeUeZdPXBLjh1Tl7NxuGmQUICuPwnMj6pkC06W
8X8UvcylYwiBcxQn7v3bZdNd5NL2d4FcyCdLesOBe45y1QE/t7hr3c20yGqHzPA8lhReVB9xEdlQ
YafO5heWRytu2WUb6bCc3QdHdCSeNYNF5qQf96KEegiVPhi9zjDaE76fddI8m8ez4HKwxIXwtUMR
iYCDL1grnAJVfeTAttUsv9RBe1lJDd3E8+BgBoti74sR5OPgb0gsaDyuKP6OQwqh5r/6e8gWJvZ3
0LCv6d2/KNjo6rffzmdwb2wiC2Fcdsx+mPy7B6nHTILuSDWfiNwQ2yjtkat1hiN0vOGk/EOltnBO
QYSTkyVUkgI/uSAcuCth2GQGzz+eXBxvYhdPQ4f86ZuuHEDjZ6/5z/77fO6BrbkSAOixpxOOtWh6
Xqmf6CAhgvtclyWmyI4UEh6KjB4Wrj9I1wpdXWf18vi7CKD4lBoUEMuKPU1V8f7z22dSVqMhlC/x
oNQZOKOpQQAtNG16sf0rVvrV9zqZkY7IdZmpGiOGnsC7GYcfqvNxFStnlbv3R+nySBmaeSUpzrOT
VbBYS7OfXpKhNlakEOKYvwnMpz7vXCLftXxpVLhCT1Ij+w4HzatjMvDkemHIwNLZDTe1fsWek8N+
NPLyup0U3xXuue+ZLOmgkWRxz1Mlbl1iTp2qIpw9/+EXljSRlhBmx9R6Tqc2ndaOaR8gIPEhrAqy
DC4l+5IyUYUaBkxgEJSwS2WO1mIGC1COwU9yRXZYcTWwADCWcToExQ6fJ5+7iIA7t1lRznps3+4J
1sSg7ao7HjI1v1ln6aQ7YQrWaxg40rKT4cY7kEEXUCuyvDFy/3mV+jeL/Nb4V+mQms+HXEzfWQ3g
ISljo7oyt0KaIED30lQKcb4rv8miG3gc+5c/b/DBjImjZP0wS8q0X3PX2nNOCoxd+rMSJOWwDQ0n
tSXtrTgn5rLvM4yiUpnBt8EoY1Tbgo6VnCvtqbkhAKzRfnViCJahY0gJS33KR2PJ62jCFT4C2k8U
ThaQ/BsYeLBRqQdTkwaUy4+uQ70GJSYT+R1su3IH9KdTeA3XbiTgFJaDyRwpORD+B4G/wZL8sotq
sogKshIV1uRpmfwXrHhUz0bF4EyPuEji9atNZ3wQZ8tsfT/5a1t5tVkJlxyEAPk5Q6GS33QR9uMi
TWRPwhouY3A+2JE0sBNrktd7q4eeaSRLja/gKOirJrjie2Hs9VOeZs+fU8eHLund0vUD7whAvzGw
ZVJkemyVFE6hgJyitRzigAQk+dC3SrQiDZCYvQ0WyzsKiFczavhep9iyj7Lm9tKjiEh7V3mAydrr
HkREBXN4l6z4UAjcfnXNzcA2rtIs3l7cmzinz8QB/QMDesAaYFBtxsYb86HRf41KsiuFgOofY5mq
BGTrTSF9tL5DeU8NIO3BrYNWJxCz1UZp51FZQVw+ZHX6LOU360ucewIb6j/PnCMzHcAtgKBkdJgI
SSSQD2RDmrpFful0DKg+fma6UVjiWWsOIFKx//jSqdrYxQgczBSF2idVOS0714naBnFlIBRP6Dsh
1JNOGeWte4zZuUHWmI3kRgnO44DLpBNrVvzBjT3grBG8VtFiKEnIbwt39BmncX/dPy0KjDsTobhn
seH4K/XlGU4hpEbMtpb+QukGhUj6Wlh7c8WpmEa1UssQWhvP3B6dzmfazJ9MSkInYxgGjEKX9KCY
QKXPbwVNl7kKIV1SaCZcwJxuNbyWegVxiRX9rcgiw6eGwF+OPPLkpOXbe2w/jGRGUp8vFkyeulNy
oETzG1cIgUxuzqi/do1f56SFFaw8NdQNyQSQa8qC5dgT2J47+J+rUwU8PGwYcL6f0geeRKKsvwZn
xce6mBiOTDABi+EYt/niPL1VGUvXQvJLa1QTOizqxXVyU2eczec4QUILEeyPTWYZEwBof5EUzI0T
OpGiDr7fMIUk9johxOPAxhWVYoBpcdA8qbYsB8EF0YlVQZ5PU7Cm7KQ5WbRTENagbYqkB2owXn1J
AmjCwXaF1XWx19SuI7HuxV3jid1nEupNvtQc7S/UbHDiHTU+PA5Wm/hAKQN0ldUU29x33kVwSKgZ
N1C/DLBEksFOr+7Aa63riWVg7/wSujWTPL7Fw/sByg3YmUkIXKs73408GwF6rsoAKdYS6WYmxMRH
7ofyKdLpEFXtUjLom1ZHpvmbrTECmE2sCk+7doS3lrWsjtEr8L2tizEn5vcAHleAREYS7yd6LKWC
hY18oaVDlsc2F/ORXy/QnC3wb/zga6AKniwdVT4iQiAsZDBjtQqtUrGvvAI7U3Ui2dlOhb4H8FRu
3Wzr82qZPW15FHDaZSIvbk2QdT/LtEjOU5GNKfZmlAuuqdMTrWVdlyLjn3SX6SziSRTSJ5K03n6U
ZcLN1la1JWNpm0tHPziwnOCVOcQK8exKD76wEZCVGxN4QvBAkpwMN6/IlY6q8SAkWSQrRXRfvwGh
tl2pT0P/48rVsc56Bbnjk/d2t50hG8EP4QvqLWiEFapf0FPNi8aubXBKS0Jl2mfcmd17nTPqUocn
jy24IpVYKQ5TQmt6oxpE4GFU5htyq9zMmdIJ5DN0uLFk/uY9kE4J1BlhCBvOlPAgRrJ0DvaZ7uWB
UpZLntNpUK6UVCnUzZRubjcQFuUotaddpGBXGgUfUSD9urwk1cN+4R2os3NQa8tA+YPFbBx8hViN
h5g1E7JC/6QO4PrhKc1uoqMdlL6r4O53/LIMDnzn5tbd6SUjCOwQvL4o9TkFD5Uy9yGw+kUQiU/F
CRgAJdaeBK+A/1B94mZ8+s/66oJcAydB1qgr90lXnKOINSAvTvw0Me8hvSYBCwv6dtMY6meKdKZ6
95CXS+wNHcaWXhxyg1rb3cG0F5JmR94GJC9PSI32BKYgGrscgW/OvgWJQGLVp5tmOgO6qJt4KWZb
lTg54W22SjX5wPjfMCez1H4jcS4JmOx2KtbnpLCrxwqZ3rpC+OM0LdLoUuoHHTk9UW4x0R52ufn5
uNS1BS6E8pJmm3dx7hP62W6EVsgNBgmG1Fg78TkZ57efNk4FuhUer0sCUEQC3Uc/sQfwUhnec5v2
pCqTj4DE8k+MepfI3HtfWWXrE0gmLSmdHRH2ggA5O+n23ZN1VeNeIznnTC5CnDABTc79GOLreMEo
NTbWNTYvMvn8F1G05+CqxNrg2Yt5hWcBjh5LO6uY8Bj4Nf98xQxLA+kXFE2K+drHQrfxU+kNi5wF
6RU6kYZf6NUttzc6cWBVGvs+NKSqlis26rlivY/SFF0flYgTr2m3GTVtQa80PM5keV/m6QSG0Ciu
JopHhF+bztVWzWb/YdDBXLAe7y3TOmmG6XvbjDz1QkgyECVdphpJHjYPqNGIuI+PwwawfzDQNoB6
/7hbf6/5Vq7UiYRkrWrnMruxr+H9zwUiOTrlRmpecp2fLFx7LDXzLcrt9SxQyvjdCYp+zHBYVTbU
yaQpRQJzuTyNlKeiQGt73EzZ47RCEoOlBJgxIUdsJwpoEUpNZ+32BVsEwCcg27hdoSGniOG9UahH
0tO7XFxjAckQf5WKnGoqRU0B4vpSM9jIl5wkrZNaC5hfF7/6ZO+sMhj2/XRwOvI5egTkJiZ4wg0P
qS6rSz//LAAplXTC/Wuty9X87oBnQGMTHiY88BpuaNMMKBJRyq2UR8d6UBUrASyMHABf/fF90J/Q
+iiAhjpRDsWrUqQGNl20W9QLK61ZT6nmIsFNwrWGajj37a1SJ9/t3cPYjOcgnXWAB3wHJotcGBMB
fFYYM4PMFPVJK2LYzhoqPPKVXJSmZE8j+l+RnbMk4f/NRgP3AFFif/Mzmwh+JV5gwxVjMyEfBmvr
O7IJDpNJndmQ4x1rL+Mg1XHNYhSuR2QSnfv081Iew1UASGneiAdlDBD2Vc8gzx6kdZLlaQIr8vOT
BiwJFrre46zq+FUjwvRCkToeL4LyAHMuxKhoECNp9wm3kAq0ezOUJnTzsBa5lTH+tCZtR5Ttg2n9
rvcD2VMFyXBbclwuiwtqR1rUKPlXYOpu1X51KrzBmKBKS2q+2ppPbkgjbJV/njsGdenHyjWfvhf5
7Hhr0WBq69cL7kz+jF+DtYdze7Ccnee3cRkCwnfuHO+lmQYDq1830EpgMTD5CPK9bJecBHwLib9s
jsmGUDzxthXbVYSlD99ENyxQLKEC41nO81xr3bghOkSRjWspcFqSSdWzAQ555q4yzumnbZr31O8f
/1WpFnBtUZIN8M9wJaxVxd11cTtOUi3Fh9jRpwa2jz/hlQuYSDDPKnXasMWJDwiAloE3l0q3WmZD
gQ8NQDoIvUP74vRq67uFcJZ4ZZXJel7EGm/ma1W0RkPJb0pKpe81d7lkOpBEXAdsXp6rYjVZunPJ
YzXO36LxJlr1wMBNbHxPEX+PDn55/5YJcocwTNTr/mgp7sjxUFvOwcf9iYeJHVL3qSq1Lu27IJQu
zA+6eIlYXXkcv9Rjy7+sELBxJ3+GbJqemFMjDZJmYcSGMQ5UK1slPlvzOHIliMcnuoAW78h2mBVj
TUS+sqUVLaxR7KjfmoHHaodZcWK5r1rA+t2Q9ZbetQEsHXexoC1IsVaqNk8+QBSqzoazNrSpLGkO
bdMD52Xs3QhXF6nzZJ3t8Gbpboxialdyy/VmJ3loaNjmm5PYvGRJR8NLpCN7QUTUZUsIXYiDauS0
GesmXSDTIqDGOfunvximJXxNRdaiv5fn+ehRUEhzDPdegQEX5qoIAonZ3tocgaF2vRJUKfdR6OUW
oM7wDmymp89rxhJ0IHoYjd9KE2hubin0Ezf4cIRU9m6S+K7rpAaQ0K/D25xcx+Y6DsQmC9k8suAd
BTJycAkybLN3eQeUmDUr4jqCY+GOZlnHFnZm4Y0snr4fVpJtbaCZojvIEM8n69ul/Ar+dLS+dBwZ
xmoplZubIk35/CaQkrhCEMJrcDtNmnTwzw4GpiyfEFqthjOuiIwWeYbg5hM+FFnDp7r7P40fwJqV
pbYSEBqu+OJIYNu80Bj+1QIfTJErnSVujh8sKatFJ02uyeN19OwkbW40wT+C+A7A8ST9b+8I/h7T
UW4Zony/tbwpFXyekuGNDv5g3SEhF0vr0Xu7Sc+wucwpQpkRa/ehOsoLPTt04SLcRUTggArwfn8k
pPWTeijPGH38AtagHJHtIED/pmn+HkmzdtnbAfjd+5M+I8mJEoml2MoObewEilq9HsrUFsKMH7x0
nXGyoV/MND8grBqtTlLG9FnKo5qgrXSfRsS4KJrW0SUcRqjRHnB5o160oau8f3V60TGkowDyZSxV
Y/YYaHipWrl/Is79gyyDxU2ofMAzLY0HHLezXASG1L+r0/BOiSDqoHFynGjsnztoVrrP7VmmWedU
gsps0VAl2h4DgjdyaFJZih+aBvT+yAMH8S5CVpGw7/ptfpxaHd9JSy0leEx4JAY72FFf+cWhYnsK
NOS7FBLfrPHKk3LQk1Tr6nU2CCMxfyL53mi+IlEcvJh+dmdCYoAeSvtV6N0CZWu3ALviQryP9xYb
HDmzYJcNDFnrVCJQOmxTJO3Dl6MIYJIczChgnEsPw5V+2uqy8Ibqkr4wkll/WyrZGSZh6TUKYYXP
8XjVVhMD63LhLzcwv/pNN8YwGZG3PRqRY8LP6UvWR7iHHGH+QmQtrX+QFUOB/l7p7eIXTvPL+uVo
CUjrVIJKcCihwhPbUxyGqtovPQmOhMTahrMfWskARJpubZTMkVIuGHhFDrP3yDTgbBhD9y6ETNoF
P/F/i8ys8eeKwm12o4/cDwQOg7rRLtUiI6B9eFjuhZkFMB6VnMknFPvOhZaJ1DqCiukdVfMobMAW
5gmXxaGHVWB/ixl9m/PRZN7/x0MH/6STNa4B9sUmp8+KQcnPwilkTozwv+sUfSSo5CLTCRry4V4I
7I3TTLrptXiGqZYzvkFpwD/QwhO9VpoYqspWHo6dvKchoTJu+73sLNgya+p8rgZD1s8VhCqE/Lda
h+cyrhebnVoiAP/2IppxJ/NelXJ/0JGiVmrgZPKgWHo6M6THWyJ8RmZvZKug82HwUAA2tfyV+ZEZ
qkreWfgDAPqoCLAsH44/h+/iwrnxJanz6D1JG6ikL5xK5GYnmTYGKOLfZBHnhY+bgV2pDcjr2S9b
8EJW9ke84PPxpY87N/cyuIMfoEnfbiS5Bf/GLZZuSAOgW9yb8XymhfkXanr1owB1Gmy/ctzaQ1XB
kaA68I7zopW5WyJ+4ajo3gs8Lhg2tjC2/TfWg433r/vs3KtS8scMeI4mAvla13+GTPG9R7JMZY4v
XbenLy0V5uoGXnpKzfFwwMFo7EfAmQkoWAJ880YwPUqj+nXfQzqPAIlMvSAsuEtrWeup96L//CER
M5XJdUJAP6/uoHgw4LkEPIBfwM+eTRyhPmnSYVI14fjVCuCbhvlPKyPWnKZHBT9G4MrK4CmvyTtK
x/F/xv0nhkA5lRaz5ZrYX+0+U9L7GuGtqNo9pabGIrUzmMFwCgdRHEIKbm/whKclXxCY1VDGEAAX
2ns0sPrtJ6cPb1ZE4C7gnK6RStLF4VGmjFMgKEmzZ6N0Ob1CoCVvT1BiZslB08YBYxWizW/WLxHg
o8iJBN98I9kXTXZmuG1EfUT3lDsdjfGsCO6Dsft8Uy8v7LsEqfssS0E+RQLAszQfytinPTX/QLOW
zdR4o9x1w5eOYcgaqwKC3AdWVmNS/A/ppjCsw1Jze1EbBuWlATQaBKU1NRiVMrQTPOzYLxmz9sRh
golBejVDMBYPGHXEFc98ywXFXBDgzdsTDGnZFNReNfe3B8e+dONToleblba5Q9vn9IcrAOfSkA/5
oBNRRpioZi8GWK3C5+/O8AboSUsuYYEqCUw4RJ/Ms88/Jhcn2XY9wzgoNHPk6WtInQT1heO+vQBy
VBOimAObtKg8e0r0YqCTgSREvrcWUJioscFYlwjh7mypx6FIOaZgnxXDrJsg+3mtIIxpjbUFG9NP
r1IxhxCJnfWtIuyoMH8GfqVp235oOzjd0cO4n3RcRrLntdr9wadgmv3Pyt/ONqYEatHr4HokC3L6
Awvukkz4kBMSIPOwIrBDMF1EImUpTq2hoNz1R+oj2YDMW3Nfz5VAtPalnXNjXEHcGAbZjYyY0Et/
mMDQ7HjP1EcVxy5yZnWnWUkb5/BrTwxuoFGG+UCRLHniRzsUGN2xaMReg2zi63lh0QEmwA3oudcc
USIqIPKXvl6Htzev2LX0kTBVTZWerm6pdTOfPRWNuQYPcExCjcWhf2W6zT2MAm6WpOR8Uv/dPxU3
5C4Zu2+U+xIkdb0yqtnpKDOMKdHDYmASzH3Sd/rNxAa9e4c+NjRbe+5yMYyiQN7XYwnXxveLrAyY
NI779+NXJ945X3/0OHSUG2f3A2boI4F0raYfqQ1+L/QNauRZEIUsrYzN23YxHwfhDLYy0fC+6mQn
4QInTebKiGTCrZ7nglQCakmx+AJJw+0me/IAuoP+WxjhoEm793PheGvYfZqOimmn1aSTyknrMb2C
JnHJuXVJ3ELUDA+yh392iCxOvJ/vt/XzU29lnHTVGQJ+cxb2ymgTHzMOoC3zzrNmTQRMLfhwbKxA
MH1tt2v6tf3dcKN33uMvBO4JxFkk26f0ZgmtL51K2IKkfosEwXY7BgJe28VbX4gSK7JoP7GXYp/j
Ao7NECzCsZo/I0u9POjjjsORYGgT9DrDrlQJ4kDwAotJQu+QotnJm/xQlk3xYT4FwC/stKUPzJQ3
Vn2pNd9UrQ+gvI5FdPHClHQyHwncrU+YQsMFHMfzBp8Dz0w+czb3AwKBq0K5idycocGKXHmxB2YX
ulaAg45peBHEwlqjZmORUqzWSRgE5V+tgm3tNu2hsH0qtLt8nBqSzlh2hHy4AsoThsB+rO7ClCPw
YjzpeTfJzf//5I5Ficy9YcJoevr89//E76IgGKSXl+grbhFR5dVHOe03VoOJVbGpUYvE0Reqt8w3
a3kjzAr4UsdsNamFvY0XaXRCvPTCvxiVYdoS9GqDDXynW8ak30sCRGjQfJ+YBYSzzLy49QUburii
9L7y+n+S/gV76QEhoP/tMDW9fM4FiD4bjpuTer9dYa0pSvGncP7ZGAvlLdvygR+gMKHJel/q3yw8
SN4JrjVDxnm7jXDF8uSQwnjD+67BEs+ZoEL7G9HtIPsZeAIUBkKhU7cblxbfusZtj0VKeiWA9KiN
nWCTZRaZZQCQH7eYKzAoVX87qdzHwUvK/AdxL1Z1dCnSefqLRUJVc0AT+mjX/koRyvcq86z4Fd9Z
FIbtQ1rpq/yBW29VrcFgJK5J+e2CuY0Dv3o9M7lj/USHBvrJiBke7RYARnT72u1AEmZDrW7+mx8R
Bx/+RWKKT9L+FVE6Ir5m8bCl0VgWxCAzfzFJ+ezl0X74sJkjgHCyBACe06ipxPo8waUB/Zfxfy7P
KlE7Y3nvt5Xmt1xoRfhmsjnVFHpZySmVlgC5EEyg/dbl9KY+2Meoubo0mf61MNCavioNqLcuHjz6
603y+/KjG2acmpRvVGRvjaYtR6tBYs1DKXu1GT/s1KtmRn3y7Fy+u5ouD6HlJxMBzzQJre3tNVU2
TJoBq8mDrLe2Dx7/cE9fkyaubwxJKxn9zTygDP8WTbRwM0A4q9oexr9vroeoXkyyxLoGmGzXGZWd
yskwr30ell4Atj2Njnu55JxlPYO0Okx2i4guR9Y35zw53lxpJ2RtRapXowyIST1R0x4Eo6meEzMK
YH5ykye69iNcMatmyRVm0ugQeGCsRramUIFuXpXIlvOlQGSDrPKGsVLLorgLxoqq8OxAi6eV9Dgp
LhVEYn6tB8Y4dJf1cpnKlilet0zTKnJfCFvs4xDa0IGf1bSR6XqoMbcdXLYFdWzDCBRFvbHJPfFK
8cIYBVIRFn0SyBxzja43s/Wuk1/KwK7NXPgGVXSHJvCSjNa6+gG20neABX9K7vVfPlCxf84Y3wgO
oXN6UDVAPBxFx2CVtk7zysNbTdKLU0Mz0CdL/ZjKZF67ESHTAN06k+ZVCpovbOVczzmycTXvrasF
inDC3Y5bllSKjf9+myVGgi5d62XIRLZTgsrezFXiIY9xsUM10LkXZQCF9Czlq7Hvj9iFpOnyfnqH
nhbpJPvoHRy8t9dDFq+sXORrR29pdg0+GAJ4Z3YLnEZcRkY3zcX6GJCEc4icyOfomlGPmbZGj/EM
arDpl15+E0VB6Jn95+jWNCLrIwL8pFN8SkRFIZvO7qn2lz796vurcqsExCidWPwLBM58h3kB/X/+
ioQTdD/oLkr5rXPfiwJQftK2iWmjPkc77lNXrbhWfRWZTID4VQoHFS0CxeqxR9hjzp+haPyXZ/y8
X3eljbFTaFu8cZjwCYQJ1tHRgyTZUzTb8ol0e1IYoQ5ItXJFjD8uGxAO9El4OYKKy8hgNXs71dEy
jAy7FThUZFErZsrDqVEvKCrcf5HhV3kE7p8oP32WN5nR1uUdgZq6mPtHtlYG9obI3frYj0JOmrzV
WZUGQ6r0EMK0cr3FLZDCay2m7+YcM7bopkyuAjRBjQU5g5qjGoECxgu7u6QFUNPzv9LmEpwmfoRE
H+wC15kJ31evVmCcBz3CmhF2AUeZw1+epnTn0lUROXEbaeZWkzlo8JCOfSspWeVL36n0FPCaqte+
c34JGu+Nd5frUMRhbjmwti6k8gMz7Wx+yxFy5gYmxSyJLWbTiEXi3kjkDJiMCJSmF5UOU+LGfM23
/T2lBCoMJk1JCOl/jZgD1VJ1adqV1Dgb6tGPhh+hiIV9t/Cfv6LiDzxM4cN/ycW8yuwN+tRdtTo4
2KoOEgP2+8Ez9hfqLojDcooprOcuh8AjyNU2Y3ckqEfEn4JOczTWgrE/9uq9EreFzq4TGk6fs8UM
0iSRMzbPqbbtgl4UVbblXQe1fvBkB7TgYhF0JcFhNlWYpm/yf58a7YNi3LZCYcikqxuNS2W1B4VI
+KKcUmkQxuDJJxXvTvBBgE2RfF+JUHPG4aV/gUJxUfvjMLlu+uxkmEcBFDOr9gGKGHsO0k8DG+V0
7Hvh9h88y9YvNAj/ZMDOI7DBCMnQO+tIwk09O6DTsFIQ6jOTwiIFA5H4tO6N9zMzZBmcFWBvW8Lj
hElMqfvtm/wSSjezFsOS5Kv75I4sYfp/kXZiSJgPdGTWyNQ/FkDh8oMnmYtjNJ+YZOviJ5YjZWQm
UKllvfqvBU2ibQ+W4la6yn9Ho5V/jCmf4uwZiuiB+HVdR8PcdeCfNNtsOmQQlkNT0QDuO4L6R24L
rGJh6igo8PWmsF6MhJTJEbrapoPBN/0LyFTT3u2qsahbcFf3hpLAD2xJcaALii0QX8iJ3xJY7Ok7
q7bbACIWYU/jYxru8o03vYDgx3A+2X4dOOE5FKFZE0LHp6l8cx456+9bQpDwXwrqX8JQbBtp2Iue
5myyfxCPzJfybb9MMfmPjyQ4GeAkusYNBdIxdz00vOYzbfddzALyUgRQ8UwuXRZ+DAMHJ4tvUg4o
ihep8w4b5lvtX1atx46aCTXjsMDh+jNatM2z2uLTeTdYowRzWQkLgHY/3Rk1rtSRBOHC8zqMOmGZ
Q3z26aMviImp1DouoS9YRk+GPBb7itJm+n1r7X2qgPXwg9zfHuOAF9oP6J5LhBQk+U4evK31eHZO
DCA8q2KDGSsZYUHbUJbT0du7XjR87lLTRXqbxq8zAzBWubt0dbNPTnYtfwSF2EeGolvLhuViItuJ
v2PrLGqb2KmtClqoKD6WbnWEQyIodN24K/kLAlBl5rUvjIIMtz70prKM52WKAuW2A6bEyw1ySqtl
KOpjTCzKlv313v4FUk/seAn6+IEPMIxjiZKvlUaM0/amJnMiNSD3/owsx8ZnbzkHzUDxPtzmA7df
ZMOrUnp7O4mtZUs1MzBmuizo8cV3xgSuDm5W/UD+syEDt5TSAFiNcnzbpajhHp+UV9wksxkb1iXi
suy3wBC7U+JNsVC1ARi2FyK+WGb1mGVuqKL5Lm6E0n6E6W+Y2dc6FDWq1csOGoXoecAF/JnClNvk
PMsOSqNd4CScMXJknNLizkkJ9JPAchiXX4JeXXoYWrLgkZEyq2KUSU1vS4SpFe9XfAzcxxEiDYpO
XtSOlpY1kmxsNTVZVtc9VcmpcRL11nDY+hcT3skprwMXgUIxCq6XLldJlJSD9y0e+YdSLnJZkZqh
1bYigu4X61NYjz1Yl4fJoq9CEIBkyj87hVtMzRNM3FkjigNr/AkYY0vTxh6HQGoI+WaRZKEZMtSR
Gt/4++beaZk0FJolScqZWTKcr9zKF8YPQmS6fs7oSUzOZskbIRjNpjzSbdkVOtiPzm7SH0LSCWf6
i6mR0dio+FWIKJ6WTZEUPwXuHSG/bgR8uGxhA4CYDkuktnmWfMusvcSDuhj2H+jBWyY0JA4RGt5G
nUFagjAi/Bc0prV6sKnzi+q9S33GCrPnITCcLJgPOKXtC1jWabEHVkBVhXnh4Uhmz159XqG5yLpD
Mh7YjMuCavqRfsr9Okdx26fmvil0H+bVqTP509m4XK1JM+bbAh93ldFIdluNwxvZwtApCu7vK859
TEVgcXGcRHZ3FPXb1q4fJZ6K+nJaJWfHFO9+FEhWEebz+gf54NqPvmGIToeeSBZ6w0hX9xpwCY3J
vQ3MHvUyMqKJxo5jyyz7sC3vYjqt4N2JvrFRH3oKLNEY27NtN2f2gdUs7O3YkKXBYK2eTkQXmRAO
THkaLWIQ9mfmR3pBb7FOFMufN/S6GFRXogE8dkPhHB4u2Uy00YW9ViaUbIKbvrfcRk8dUACQEb0v
gffEVMwwhitWCGId1s1kcCD91lhJuOZYa4mLYyVimp+0wN8oB4ISEaPhVymnQysTpqfSdKD/LXm4
p1qHUi0Y/Oj6KYiA64QV86Be76XKDfb/mSZxyruwXT4QsOKfnknTrN4MfPTaZBj6UW1h95z4Wl+9
XGAhOJ1VsbyluN7hoADBS6vfMCW5I2NSsV4hXP4XulRIf7L1z/VVyCI06SBB1TkfiuqeeGLYscfz
Df4BKCLXNxcFCHz7KuxUVMT0xLvUXtUOJdO3TaFQTBT6OrTq/pTcZFW4ky/HcT60dodow4LbkgFQ
hE7n/O4WCcY2uUkszyMZyLjyhnqaHRw51L8MNLPc5k5lzyklV+72bwguDjdJC6PbV8efZHkQUSwz
zGzUnpeP1LCd3edtdz2wNkwVcTDmOpImSsqexS/niHPNPoGWJ+6U23MZGYpKMcxITzcdvZrbEwRz
kw1CsggDTtXjAxiflu4d0FHp2Nl8akQ37wFFdqYIejUmuurptIi2rOhEJkp+wxtW2nVbcq41mWMN
Nqi2CfPK55hPR3ZDvIpAPs+2j0Yi4cQb4GlvKuwNR8p02P4kixL1JY+sAEIvs0xezMsshUW0H3i+
l7gI2YrSMlbBBn+HJHGwdAScnpTUZ/8iPb8ynZpbRLO+aN8UmWlb5bGw94sG0tnsd2nTl42T579A
JvgUCOlMx566D8Q5cO4P3kHbSpH5BGoxD1io20hgGmhq2Cnv38FxvmEZ9zp2H3NY2S3wCQvVZtu5
OFYHE69O3I2aLDPBu0+N6G24R+nbBJFxKTQ+0BZLT/EtnAb6kjNnmJRrDXc9xdPuHO+lJgIK7JJT
z5rkRAUT6yGV9VPL/NuMmvih15H/weKm9/D9GvteSGHsQgrdeyDBGbEeHAWlIhfDns9f9l2fIn2e
fQqs6r9y4/Kneff27yxqllS+kDF/vVRso60nujjYjmxbDSjIRo5JIBL4IqtpbfqlVq3RmvNH+2mP
a21e6CEWBfJ2zMihA3uhD8l36elcj7V1E/mtPzpZh5i5NNgQtNz1beCnl3OM27ppU0qwghoN7eAj
FVLEVuw25yMYIKi68dXAFqhl9cR+UvdXlU6JHVR1bvKm9EDlNSUrM8Tg2z4+hbnk2+AVuDcHaKSA
pqgh5CLY1pJzLyOytzVbwXTbqs/+0ZZP1tVUbt9UTslhc6RurBVJJD1P57RfSHvZv9bLaAmgGl4e
OjlI0paWdv2KU9GqtTYEV9etA1oOc4e4YdB83UWW2W1HC9itg2O4QH+5EVwsR5yFHy36FSrRF933
MjC6doqMS5IRsT19itoaNjXwth/yOF2HFed4YNrwFhaNeQkU9qSfa5wgiIzwHZDKV7wTozlx2YCh
h6C2U7aug2m3k8TCuCFEzJ4pWAwju0HjOP8/Ea34ln8OgvRnH7sI52pSdN5NAWtNBbP7dYoOELPe
JeNdd5G7q8/lXzD18Ux+HIWsc69YZEXDi327/+i+OpvYzSg0q3aRjQvdptPpljuDVmiBy/XRSl13
PdxsKgziIMW9KvZsOxpR2zjPFmdGuPeO5JcIi/Xas8xJoeyKKPkX4YhMEz5VXB5rGqox6HWy2km8
4KqjzBJmxbHiVHT3pgVnYnq1P7QwCmpbjEFDKseWZifUjjIm+u2qjQG1DLqkZDsPpfTwC+WwoAkf
H7eE0tL0pyjNJUh8R9c7rdVMY59VY3TvgMuSMvNW7u7hOsLp2Txtm3PpRIiuf/FmCIggKH4WEB0/
d/QtlNEZxCLBEUvmvEWuo2kgNvTJiHdd3RmwXvN4zbyMr4kmeZjZ1uQ5IJqj7ISq8/htJqxGfVse
5hrRYpeMIWcPPHoM4mY2Fcgm5Vx2Z0bMQrVrs4K6u1+6ZrGvbdy3Z88xtXLYa4N9+zdY/vmEG98F
pZltnsEo9vfgGC8pUhySiBfw9zGj2i/YFKVjiME6h8zy+MQvc33ittPEGyRFzugI95S/vpCQhscJ
QYSlJSp0SFG+TMNUDSremKHakNK6yEKsbQbSslOxHs+wgUH+oGj/OFWKcDoACaKdTAKjZFVec+na
oLtpLaNsZkeJ+DRchdgodAkDiEveTuPJjtXKXtjH7KUmxpXtcgtmSRKbvNSvZKH4BRPMX5x52zQ4
WJJhUBCEWKoK9XLdeeVc3VtU1rsk5UiOyXmUE4ssbE3ZDcY7WxZzDJe0/slOyiwqX+h9N3NdGloM
QZA0+kr9cTCe7YUeY/H6z6k2BP1t7pJifNS0xF9dxRBnYGcct9iYm2Y9N7aP3mQDVq0qZ3pMFsjO
M1j1x9euUyRjjIWKTI4SeZ7yp1GDl8O5AvgLjikOGwj3IaYPeQooZ5w7KDIrrFw9fgIb4sEadpiO
UXtTGYTlzqpeqNOPvUzOs2+XaMFaBKNRS9J19OiAMxuBJpDvCx8+4AY2okLcel3Ttw965cz0OSo7
P+aTkoml9YvE4WZgJDpxpHxCUPfa2qfQ/NRRYOAOkw42+PbB3wRtz/snMzuM5eq5P5JzqJ5z/7W/
+EPzW4iN8wWoRvwE3oZgs8v4NwmqeEjmxjPBVn/D9OUyXGPt6ldnpDye/ozen+gDGpjmpOzQofzj
1ZfB0JYp2ZBjkU+CtQLf5UPD0ZKRe+3YhFgbPJq9tyJpUt08YLR4aV5kfxKIIeEG03w2xRiIo00d
CdS3d9s7Iycdh+xQOdTtBsKPy9mcB8a26HEUgrfPubgTcZF3s0RpyAp0x/Ul4ob+bTXm1pQuxMm2
R9x5UoeveqIDFb8a/In3XbqfLjqHmz2HU0cA9JzZC8JLu4ncCLjuo78WHe/0rLIfPKSCFpYdM7GM
jhv9m7Ilq5+eNptSL4CLGgsZLJg5YnlQcQs5XJl2CfJBp1IFkB0LV+q0/s9BXOGHyuV4gkdbL1Ok
RfAuKVs3+wvBZuubJGtQsQhZphu6SVzdTwrJd9AfInhv/pyR3mrUnrUuIS+IBG4st69rTEgx6NDp
UE1msbcOHtj1A2RQ4HP+jI7DxgmAOtKwdh7BCQIhtl29YoBTIh+o0fCS0N0IK39syDjFIjRfo+ro
OgvjjxIXGEfTGdk83TQ0HEZnDnUZpQhaC/x0DL8CF4Cw7njf+l7kKPZ1i2xNSFOMB9ud1II8Z2gz
sK0hjZlQwErBGpQ1IiYzMath5NgtZY1USZHFnK9+LfNibrwP1MVQHpecPmM7VMqcoVjtCdhfa0I7
qmHAaWLrNImTW7amV3hB33yWP+5UznKHpQW69YdnDBwUEn23WZjPqtXP53JeCSNrLITSVGPpEv5L
5GUqdQ9GfRQh7b15zUw+E6X7Y2N0Zkg9bVEV3+LUnvWrj2U95rVzeK+t33flymjfC3JofPKGq+q/
25dZHkjsxbAKQ04EW8Q7M81TIClVkmVD20jteaRZtbXz4YhAfdVp20NT+pTkmGq9kUZv7mEOEi+g
97dvmcWIajUgmejchI4EFgmR5gXkA/E/lkyl+sNTW+pi2TuPRRhKpI/1mcnIC2g7Gr8xfk0mEdKe
Pn9bjsiCvH6SKIz8tiRjBH2FMieW503fQy76tOIDn6FROQvMjh5xROqqAjO31ohDcUCelKy3llTX
2f5CKDFF1BaNnk8Pw1eLJVgibeN+tfKFv8EjHEpPUhCCj4FN1yqgKNm5B99VF2cpAzqN7cC4rX1C
2ABHg1M+O87X3xFKcXnGNy9tlAtHMd7PeNUb0ybSQ4JJnNrNbXxuipYgdiTX53ApR9iyMNt0jn8Y
tUjpRs0UGF1frdbAPBkh6sIarK6udu1PMVYE4rHmqzu52WSAcGgXM7Tpg1iBtwgmDTi3FWFH1nKr
usdeNA98RFmdr8hoytmJq2K52I5pvh/NSiyJYw+Z6jjey3Qzf1DW3IaD9pqWTFFhH5inxDRKqJHX
/tyhag/D8IH9N8BMgzli0obCPyj/v3Yj8LTBl47AkztU8znwOfH9JaXnLmgZJBPrKESB84SIXUBW
ebEDShhuaPupvO69TNV+q3PlnV2BtYfVL+cityvShDLvhEKubtlV9mPIXEQQ7tkoyDy/W8fudXQV
jA2KaivSiOgyqsJbAWUPl1eYgLxLaxEsHb4A9UyyDY8IJMm8yiq10osEX1p9LW97LCkD1RntMKVP
maP5Frs6a6aVvICjlgMpyyhm66ZmEyUd/2MnfS477TPaIxIKTQmiNza2dmf9cuXM98c8fFhOFtVs
Xywls3G1eIcP7DVOBGe8iG2zk3+kzHCPYznoQoZ9jm4m8Tx0hz5qoI1i8Xe2c6Sfh5FU7KsBzLMZ
Kp/58/iaVCp5PoIpaB0u7SXLGIeUBbJANvuREEmJj45Oc2mnsvIA12IIKX9tOAcMwZ3K5TXwMH9Q
dxULGQ1IhPikffAyczCPSi1z6h1Nv2DbkD+FThRZEo64DH32B/O5I+6RX28Mj57+VjS6EtXAYBb6
OjtapgWFQqeX0xnN9LSaSrNTzn/KJDC7N0uGkWJZjNxqI0Lmv0MGbPPO2EWqG0EhWiBZlxaKQcRw
yi36aZIVpSw3OR8ptdZKdehpYHypOMiRaN6x0DFylWOTvht9MOyWs8cIalRNhSgRkiHUTqOGQt2L
c18sRuts77cLRnsriwGkfdlR7m7mF2IuuhLK9D9bxx8sb/MKLfM/nNtHMlPamHwWK4W8pZDbpj57
F3nAiviKfFWTenrsLW1CPQ9fR4j/vZ9a06HdWItbUyYeFqmvZGYqRvNDeWvR8m259TDHKzDu2LxG
5S3hrptTEug5wFKcNwFE1sMnma1APNIG9uWkn/G+Hqb1Z8YtieKz3E4YnUPPJPZ2ilf4gzjxH5jl
/FEOR4ixFZ5OAZa+KOemesjUV3beMbYTdEVx4gVFTGBs2pNNzJo9f9TGci4i5qWcEAq5cBiCfmX9
iEyIlHJQaKe3oQUBZMWlsxUVckae3GOvXQRDEcFc+CrfLILjH0DHAjFqQryzpng/gBy2YtV+RyTe
CxmGZWh2Iq6HfjxuDSS7AkvGAv2EElCOg1VD8fLtDtTd02dAcPF6zq4tBAtPlFbjZOZgJPY2Cu9z
bc/anzZEIHkrpvOetl6dxVTrzcM4vTJsR3a5YbWtEzJLVPZMrVUzYdw50RhR/AZZ73bhXEvEpN3X
bk0xmDZaa7yIcoc5kjZzxJtCN8tjROKbyV4R8eO2Ea1VrqD9REGXxJFNxGWp5QZPY8/tJJC82H6W
PXAtt9mClxZILS81exsq/5gQ6o5mN4n3b7UPOyLJ51PCdBS71G5gUgVvjUp6/rcIsLjefCBQvuF1
QcZvd9zHc6+EUP9Iet2vyVhs+sfqGBHBzyWVwGVOr6IEF4c9yhhQzSXeoulSoSXb01juK7Z1tkC8
XkSC0AMqG5jkMOa4ovFufYyKP1SGvYA4iuidlgx48TyzHn6QhaRbYu9MuiEJKa4C6mJ+llaf8GCH
GKPV01/AHfS9xNzae+3+9dMgpcfv57j9ffVvx1s9iqbT4dlLduGTe4GClk3h2SB65JoP1WTx9nUc
44USg9c6YFVVkbXQR/y8X1I3h8sPQeO8eXJzK6ej7ZwgFuYqwxFDqPq6LALsoAsjL6d99RzIBFbb
cVxGM29SLtyOW3nvjkrb918nh9yDP7fFS2lbb4RuVKHN/AxMbF9ov23ncBHCy4n2lVPLgdOx20aj
WaYWXEPlGQf2z994/MelFivCHj1w/xK7jq1xnuo3pxQAyNI1E/IMRw6ZzxZ2C6YLtN1jluch4ZcT
iVxu7+TtXTtGobhpA+dFJcjc6gHISRJYKXMF4HNZeu4R0D2bJY1E081lMdv93z4IPQ/NF1OhPXli
sOvPs88WbIOQvF8Pfw7NMZOFftDW571vCVwCaU8bNywisCS0zc7bTLEQNtoADS1QoJCpi58hjiwf
kZPtMLDJvZcHv3dYTEn4uqOv8T1g+/cY2PCTvAGyBQZSjuqp4RoNdbHhH2wYjF6zKJYmxZC3fMH+
FAin2Ie8R1XTsxANHt3tE+jfB1UaouXDMXFPCgu5qlUAC4JV+7aJmDij+L+B+TnlpwUCFoXSreCd
bsv1H4tGRNESSdJjCD+V25s8qjSo4IwxaQOFT87LlRGTf5HiSG7X+LathJyhl7yx2DbJL8/NzsPn
mR5yLtDX7rabQjVgIRUGsoKcS2JKi9zlr1IIrUSc3KwrnMLIy2dH0e+dWJAyyK9kfbh2UIROd5JM
q32M1OsKUcOL6L21JoEhL4Hh+WSwLJ0B+b+OAGz7u+Xo19eEnALG2VgBzUWii30cuPg0yZGl47Ia
ITiisjy1qJIxKdJw+yfrDl45NVbBpzfLkEiwLFeB6YMqjhIFaXy4MilIJQ7AWSYY/Tfq5Zp7BEG2
Wpy9JWvjwx6pnccI5QdGOMafI0tZOvOiwuYVlQ1FqixXLlck2WBmVCCHCk1PZlrkuCw5K5PrtOZL
i7ESMOj+YxQ+csoiyVJWKJ/MMaLhjDgduaGEEYJwQFLQdpxW/P7vkg/RX4jK/+3XtLFcFmSFdfHR
iOPDYzN3I3ljCBj3NjCHWyuhGx5X6eThC0YO5X41+snxcjtzrsA+23KMsAIN6vX7L1e+u11iYztN
6HfzroaqcQFcsWxiO2lgn0Uxxi2O6OigNflDhUxph+ecCL9K37nF+nN9fXY1Q8LvX9ycPkqa+EgE
RBU8xkGcgmwo/rgMS+jziix9hi+BZfUAQ9eAJoOXIliBj9u1xR4Lf9ezo0e3e029lKkZx0olb3R5
nNm6yWHVq6rUoOqIFaTGhTUW+PE+ta/eTjRYKrG3e7ZUmIM/TRHg4hY49pLwfO+vMW3owryzFU9s
AI+nxzqJTR1ds51PdTZOsSTbz1af6OdV3hcsZTj9FNhPmKwuaou62AACvBtPo3HWsNGAjpgqjJw1
pI0OzU8G6Xm9EppsmFi59gfjii+BNB5zaciqIHYRzxLuEdqrcPzRhyhEYsX7TET56MvtF7NTUPln
yV3E3f061atXPB1tp5xpUEeo70y+wyQROl4x4EpvizJ7c1MiY0KEp9RoDFvlhR2hduQ2Km69RlJO
MXxW3nKUkMoL04uX+czHEPczRbjVLSjpUGXDL3/sVtcl+jfaNdIB7EQyHF00scO0aCa6FdfgULqB
KPr3Ila+ud65+YaiWx2EfSCVsh8FZJx+7Qbsd6j/RV8S3l6DVjJeuc+YO8riQBFQ7pWbBC5lkvaj
tU2psQ60HP6sNwrLtplheEYHvsRzqxH2QhFLFY4xaqliDXGzxbt9PjvcCB0HWrlI4pzw327501It
Es8+ZsTVrPlnwSwPtXwS6f6b8H19Ubo7JupKznZtAk2jpXU9K9ibsV9StWj+sT917NhJjon6QJkF
ZE4bwNQMp7po7cydHwsxHAZ/2yjOqCeC019EHTv3o/L3Wq9jobSEMrIQqUY5yNOBEQ8TpBwPhA3W
OiO5tgq6I/S2wxeNnyAceD6YUxKVBDzbT6VTvLldZfxnrI27pVpARNTSrxBUiceRTOeyx+Q2mQjz
SkEOuYTM9QsZkNXLbwt6Z1UytjXosXrZGmZ5egQkSJ2Vqc7FN3xxdM35X/HvSHiPz3XXo6PZ43yO
GpI65rtzzmOPzCW9KKdnTeWkdt7M4hkA//1OXoRAdqdoHef3Ca7ftKgxIkpJ6UZ8suRIHdV4A1Ox
vfoG1axtLjEU6rIc3kYb9kyAk9JM+xDzpWJTEstTaa8WMVPCiMxnqEWeu47/Q48pQ1Ebo+9NtuTP
+xWUpD6I0HoWlX589qvXhC+yzX59Y9C84l0fS88ny2tnBQ9pMVjh2QdZ7JQxyovYrnr1VoIsjcGw
nQk2wpJL0r0dcIoLp19TBvlJh2JNGki250AJJe6ycpDWU81rc/H2O+b/Yd/UcBHqljuUO/XRP0SH
6B8wYYNmzZ3A8yHrqpFm+u8KEQ4bpq0YGGnt1xIjpRp6kenrhvHLBO6nYHq4WAyhuYBbFCPZSC90
qIlzTOVo8a6VsUcjdCnq2IbcA1/KNyPKFrJaR7I8UPYUso1GqLlZlwCemT08wCejWATWbqrDiNhH
K7EArcSL/TDOUyXIZrp9g2a9ToBEvA6Iu7TBbhEdqkgjfN+bGOOyfHngRu73nIL7S0Aa1jE7F8ay
ZU8fkca5csEoHLhCX+lAACp1ZJkHvycC9eCxPFqclety3t8maPtHGoR3nhF1WuSkq2T/WBnR/xny
BB6G73sNrz5kxKAYA7ROSbDTqQ7a9UoHXGvbEQMWaW5IYNZrOAJSTeUizHAKDBsMgK/d3AS9B1TJ
JB1hmz64Ib3SbGzqkK2DTOFqoMT3+w0BZxWpUzCS0gJhcik/092hWm2UGsULbojyFKA7IysvLm91
HNNtw02yxyt6mfL60BCeM9waZA6CiguaIuKTXjNt1oZvaFQkEJ346MXxitfvwxsuqEX8V+UP28gM
ZMoREZky5vdRGJChTQUSC5xcCW+hsb0dkkAQajQzMdBclXSD9f5qyjkqsi/ngXLXvVbr9XZCZuNB
dLAJcpMh57lyj1OGWf1GSqejqBv/4bhTdWOACT50rOrOu5AXSLxBHp2jGfIFxOhjJvlT8Z7oxsI1
6Suw0JfpNTOZ1qWxUNLkiLsqAZaFFHtTtf8+FqzsX0JAxalonb4P6Lhx0ysd+dQTDGkK8kSXt4c3
hcGzlar4W9RxwIia6Alk9VrCdHB/h8DSQgVV8osqp6bfFtCzqCaCynZjosOPzMB7hQUTqFM5jgDE
PlTNwbW289Wlp8ZuYJcsPdysPuoOfgBA0AIRrDGwVVNLAvVfeUrBiAqkwtqHzathmRLxTBVPQvOG
mCYu7wRWtmafH3lsDnrgBv9hjxGrhAVAmaKGkHIOoD/Vt9r9HvIxJIq2Dm20iYDypBa+JwbUWszS
pLEW89/19igeKjz+qt4894RljM/I9cmrfzr4uD3b4XzzFQxAeBzvKGWyMbjc6LwEkE4SKxTMCs2Q
FGZgbOPie1qhDO24L6Jnl27vVilBpX1Clfutruo0MfZP5w==
`protect end_protected
